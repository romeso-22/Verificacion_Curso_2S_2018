module binario_bcd(bin,bcd);
  
  	input [3:0] bin;
  	output reg [7:0] bcd;

  assign bcd=(bin==4'b0000)? 8'b00000000:
    (bin==4'b0001) ? 8'b00000001:
    (bin==4'b0010) ? 8'b00000010:
    (bin==4'b0011) ? 8'b00000011:
    (bin==4'b0100) ? 8'b00000100:
    (bin==4'b0101) ? 8'b00000101:
    (bin==4'b0110) ? 8'b00000110:
    (bin==4'b0111) ? 8'b00000111:
    (bin==4'b1000) ? 8'b00001000:
    (bin==4'b1001) ? 8'b00001001:
    (bin==4'b1010) ? 8'b00010000:
    (bin==4'b1011) ? 8'b00010001:
    (bin==4'b1100) ? 8'b00010010:
    (bin==4'b1101) ? 8'b00010011:
    (bin==4'b1110) ? 8'b00010100:
    (bin==4'b1111) ? 8'b00010101:8'b0000000;  
                
endmodule